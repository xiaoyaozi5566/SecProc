//========================================================================
// Memory Request/Response Network
//========================================================================

`ifndef PLAB5_MCORE_MEM_NET_V
`define PLAB5_MCORE_MEM_NET_V

`include "vc-mem-msgs.v"
`include "vc-net-msgs.v"
`include "plab5-mcore-mem-net-adapters.v"
`include "plab4-net-RingNetBase.v"

module plab5_mcore_MemNet
#(
  parameter p_mem_opaque_nbits  = 8,
  parameter p_mem_addr_nbits    = 32,
  parameter p_mem_data_nbits    = 32,

  parameter p_num_ports         = 4,

  parameter p_single_bank       = 0,

  parameter o = p_mem_opaque_nbits,
  parameter a = p_mem_addr_nbits,
  parameter d = p_mem_data_nbits,

  parameter c_net_srcdest_nbits = $clog2(p_num_ports),
  parameter c_net_opaque_nbits  = 4,

  parameter ns = c_net_srcdest_nbits,
  parameter no = c_net_opaque_nbits,

  parameter c_req_nbits   = `VC_MEM_REQ_MSG_NBITS(o,a,d),
  parameter c_resp_nbits  = `VC_MEM_RESP_MSG_NBITS(o,d),

  parameter rq = c_req_nbits,
  parameter rs = c_resp_nbits,

  parameter c_req_net_msg_nbits   = `VC_NET_MSG_NBITS(rq,no,ns),
  parameter c_resp_net_msg_nbits  = `VC_NET_MSG_NBITS(rs,no,ns),

  parameter nrq = c_req_net_msg_nbits,
  parameter nrs = c_resp_net_msg_nbits

)
(

  input                         clk,
  input                         reset,

  input   [rq*p_num_ports-1:0] req_in_msg,
  input   [p_num_ports-1:0]    req_in_val,
  output  [p_num_ports-1:0]    req_in_rdy,

  output  [rs*p_num_ports-1:0] resp_out_msg,
  output  [p_num_ports-1:0]    resp_out_val,
  input   [p_num_ports-1:0]    resp_out_rdy,

  output  [rq*p_num_ports-1:0] req_out_msg,
  output  [p_num_ports-1:0]    req_out_val,
  input   [p_num_ports-1:0]    req_out_rdy,

  input   [rs*p_num_ports-1:0] resp_in_msg,
  input   [p_num_ports-1:0]    resp_in_val,
  output  [p_num_ports-1:0]    resp_in_rdy

);

  wire [nrq*p_num_ports-1:0] req_net_in_msg;
  wire [nrq*p_num_ports-1:0] req_net_out_msg;
  wire [nrs*p_num_ports-1:0] resp_net_in_msg;
  wire [nrs*p_num_ports-1:0] resp_net_out_msg;

  genvar i;

  generate
    for ( i = 0; i < p_num_ports; i = i + 1 ) begin: ADAPTERS

      // proc req mem msg to net msg adapter

      plab5_mcore_MemReqMsgToNetMsg
      #(
        .p_net_src            (i),
        .p_num_ports          (p_num_ports),

        .p_mem_opaque_nbits   (p_mem_opaque_nbits),
        .p_mem_addr_nbits     (p_mem_addr_nbits),
        .p_mem_data_nbits     (p_mem_data_nbits),

        .p_net_opaque_nbits   (c_net_opaque_nbits),
        .p_net_srcdest_nbits  (c_net_srcdest_nbits),

        .p_single_bank        (p_single_bank)
      )
      proc_mem_msg_to_net_msg
      (
        .mem_msg (req_in_msg[`VC_PORT_PICK_FIELD(rq,i)]),
        .net_msg (req_net_in_msg[`VC_PORT_PICK_FIELD(nrq,i)])
      );

      // extract the cache req mem msg from net msg payload

      vc_NetMsgUnpack #(rq,no,ns) req_net_msg_unpack
      (
        .msg      (req_net_out_msg[`VC_PORT_PICK_FIELD(nrq,i)]),
        .payload  (req_out_msg[`VC_PORT_PICK_FIELD(rq,i)])
      );

      // cache resp mem msg to net msg adapter

      plab5_mcore_MemRespMsgToNetMsg
      #(
        .p_net_src            (i),
        .p_num_ports          (p_num_ports),

        .p_mem_opaque_nbits   (p_mem_opaque_nbits),
        .p_mem_data_nbits     (p_mem_data_nbits),

        .p_net_opaque_nbits   (c_net_opaque_nbits),
        .p_net_srcdest_nbits  (c_net_srcdest_nbits)
      )
      cache_mem_msg_to_net_msg
      (
        .mem_msg (resp_in_msg[`VC_PORT_PICK_FIELD(rs,i)]),
        .net_msg (resp_net_in_msg[`VC_PORT_PICK_FIELD(nrs,i)])
      );

      // extract the proc resp mem msg from net msg payload

      vc_NetMsgUnpack #(rs,no,ns) resp_net_msg_unpack
      (
        .msg      (resp_net_out_msg[`VC_PORT_PICK_FIELD(nrs,i)]),
        .payload  (resp_out_msg[`VC_PORT_PICK_FIELD(rs,i)])
      );

    end
  endgenerate

  // request network

  `define PLAB4_NET_NUM_PORTS_4

  wire [p_num_ports-1:0] req_net_in_val;
  wire [p_num_ports-1:0] req_net_out_rdy;
  wire [p_num_ports-1:0] resp_net_in_val;
  wire [p_num_ports-1:0] resp_net_out_rdy;

  // for single bank mode, the cache side of things are padded to 0 other
  // than cache/mem 0

  assign req_net_in_val   = req_in_val;
  assign req_net_out_rdy  = p_single_bank ? { 32'h0, req_out_rdy[0] } :
                                            req_out_rdy;

  assign resp_net_in_val  = p_single_bank ? { 32'h0, resp_in_val[0] } :
                                            resp_in_val;
  assign resp_net_out_rdy = resp_out_rdy;

  plab4_net_RingNetBase #(rq,no,ns,4) req_net
  (
    .clk      (clk),
    .reset    (reset),

    .in_val   (req_net_in_val),
    .in_rdy   (req_in_rdy),
    .in_msg   (req_net_in_msg),

    .out_val  (req_out_val),
    .out_rdy  (req_net_out_rdy),
    .out_msg  (req_net_out_msg)
  );

  // response network

  plab4_net_RingNetBase #(rs,no,ns,4) resp_net
  (
    .clk      (clk),
    .reset    (reset),

    .in_val   (resp_net_in_val),
    .in_rdy   (resp_in_rdy),
    .in_msg   (resp_net_in_msg),

    .out_val  (resp_out_val),
    .out_rdy  (resp_net_out_rdy),
    .out_msg  (resp_net_out_msg)
  );



endmodule

`endif /* PLAB5_MCORE_MEM_NET_V */
